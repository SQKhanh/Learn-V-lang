module model

import khanhdz

pub fn human_gay_oo() {
	println('Gáy o o gâu gâu nè ? ?')
}
 