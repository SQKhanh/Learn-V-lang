module main

import khanhdz.model
import khanhdz.animal
import khanhdz

fn main() {
	khanhdz.concac()

	model.human_gay_oo()

	animal.dog_sua_gau_gau()
}
