module main

import khanhdz.lua
import khanhdz.model
import khanhdz.animal
import khanhdz as khanh

fn main() {
	println('Start')

	khanh.concac()

	model.human_gay_oo(123)

	animal.dog_sua_gau_gau()

	lua.print_hello_from_lua()
}
