module animal


pub fn dog_sua_gau_gau() {
	println('Sủa gâu gâu nè ? ?')
}