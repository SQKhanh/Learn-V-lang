module model

pub fn human_gay_oo(a int) {
	println('Gáy o o gâu gâu nè ? ?' + a.str())
}
