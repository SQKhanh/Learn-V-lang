module khanhdz

import model

pub fn concac() {
	model.human_gay_oo(123)
}
